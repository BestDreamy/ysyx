module axi (
    
);

endmodule
