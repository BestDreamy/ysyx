module axi_Xbar (
);

endmodule