module axi (

);

endmodule
