`define ITRACE