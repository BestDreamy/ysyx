module clint (
    
);

endmodule