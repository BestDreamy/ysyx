module seg (
    // convert 4'bxxxx to a digital tube
    input  wire[3: 0] bcd_i,
    output wire[6: 0] hex_o
);
    assign hex_o = ({7{bcd_i == 4'b0000}} & 7'b1000000) |
                   ({7{bcd_i == 4'b0001}} & 7'b1111001) |
                   ({7{bcd_i == 4'b0010}} & 7'b0100100) |
                   ({7{bcd_i == 4'b0011}} & 7'b0110000) |
                   ({7{bcd_i == 4'b0100}} & 7'b0011001) |
                   ({7{bcd_i == 4'b0101}} & 7'b0010010) |
                   ({7{bcd_i == 4'b0110}} & 7'b0000010) |
                   ({7{bcd_i == 4'b0111}} & 7'b1111000) |
                   ({7{bcd_i == 4'b1000}} & 7'b0000000) |
                   ({7{bcd_i == 4'b1001}} & 7'b0010000) |
                   ({7{bcd_i == 4'b1010}} & 7'b0001000) |
                   ({7{bcd_i == 4'b1011}} & 7'b0000011) |
                   ({7{bcd_i == 4'b1100}} & 7'b1000110) |
                   ({7{bcd_i == 4'b1101}} & 7'b0100001) |
                   ({7{bcd_i == 4'b1110}} & 7'b0000110) |
                   ({7{bcd_i == 4'b1111}} & 7'b0001110);
endmodule
