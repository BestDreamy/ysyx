module icn (
    input clk_i,
    input rst_i,
    axi_if.Master axi_mst,
    rv_if.Slave rv_slv
);

endmodule