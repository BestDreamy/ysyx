module csr (

);

endmodule