module axi2rv (

);

endmodule