`define ITRACE 1