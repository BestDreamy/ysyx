module icn (
    input clk_i,
    input rst_i,
    input axi_mst,
    input rv_slv
);

endmodule