`ifndef AXI_TYPEDEFS_H
`define AXI_TYPEDEFS_H

typedef logic[3: 0] axi_id_t;
typedef logic[2: 0] axi_size_t;
typedef logic[7: 0] axi_len_t;
typedef logic[1: 0] axi_burst_t;
typedef logic[1: 0] axi_resp_t;

`endif

